module codingClubIndia;
    initial begin
        $display ("Hello World!");
        $finish;
    end
endmodule
